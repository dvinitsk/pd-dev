// ----  Probes  ----
`define PROBE_ASSIGN_XOR_OP1 assign_xor_op1
`define PROBE_ASSIGN_XOR_OP2 assign_xor_op2
`define PROBE_ASSIGN_XOR_RES assign_xor_res

// Define other probes as required....
`define PROBE_ALU_OP1 alu_op1   
`define PROBE_ALU_OP2 alu_op2
`define PROBE_ALU_RES alu_res   
`define PROBE_ALU_SEL alu_sel    

`define PROBE_REG_IN  reg_in
`define PROBE_REG_OUT reg_out 

`define PROBE_TSP_OP1 tsp_op1 
`define PROBE_TSP_OP2 tsp_op2
`define PROBE_TSP_RES tsp_res
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd0
// ----  Top module  ----
