// ----  Probes  ----
`define PROBE_ADDR        pc 
`define PROBE_DATA_IN     data_in
`define PROBE_DATA_OUT    data_out  
`define PROBE_READ_EN     read_en 
`define PROBE_WRITE_EN    write_en 

`define PROBE_F_PC        pc
`define PROBE_F_INSN      insn
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd1
// ----  Top module  ----
