// ----  Probes  ----
`define PROBE_F_PC pc
`define PROBE_F_INSN insn

`define PROBE_D_PC        pc_decode 
`define PROBE_D_OPCODE    opcode 
`define PROBE_D_RD        rd
`define PROBE_D_FUNCT3    funct3
`define PROBE_D_RS1       rs1 
`define PROBE_D_RS2       rs2 
`define PROBE_D_FUNCT7    funct7 
`define PROBE_D_IMM       imm 
`define PROBE_D_SHAMT     shamt 
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd2
// ----  Top module  ----
