// ----  Probes  ----
`define PROBE_F_PC pc
`define PROBE_F_INSN insn

//`define PROBE_D_PC // ??
//`define PROBE_D_OPCODE // ??
//`define PROBE_D_RD // ??
//`define PROBE_D_FUNCT3 // ??
//`define PROBE_D_RS1 // ??
//`define PROBE_D_RS2 // ??
//`define PROBE_D_FUNCT7 // ??
//`define PROBE_D_IMM // ??
//`define PROBE_D_SHAMT // ??
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd2
// ----  Top module  ----
